`include"./cross.v"
`include "./dadda_10.v"
`include"./FA.v"
`include"./HA.v"
`timescale 1ns/10ps
module geofence (clk,reset,X,Y,is_inside,valid);
input clk,reset;
input [9:0]X,Y;
output reg is_inside,valid;
parameter S0=5'd0,S1=5'd1,S2=5'd2,S3=5'd3,S4=5'd4,S5=5'd5,S6=5'd6,S7=5'd7;
reg [9:0] nTx,nTy,nAx,nAy,nBx,nBy,nCx,nCy,nDx,nDy,nEx,nEy,nFx,nFy;
reg [9:0]Tx,Ty,Ax,Ay,Bx,By,Cx,Cy,Dx,Dy,Ex,Ey,Fx,Fy;
reg [4:0]state,next_state;
reg [5:0]number,nnumber;
wire n_valid,n_inside;
assign n_valid=(state==5'd24);
assign n_inside=(&number==1);
reg [9:0]Xx,Xy,Yx,Yy,TAx,TAy,TBx,TBy;
wire IO;
Cross EF(Xx,Xy,Yx,Yy,TAx,TAy,TBx,TBy,IO);
always@(posedge clk or posedge reset)
	if(reset)begin// asynchronous
	state<=S0;
	Tx<=10'd0;
	Ty<=10'd0;
	Ax<=10'd0;
	Ay<=10'd0;
	Bx<=10'd0;
	By<=10'd0;
	Cx<=10'd0;
	Cy<=10'd0;
	Dx<=10'd0;
	Dy<=10'd0;
	Ex<=10'd0;
	Ey<=10'd0;
	Fx<=10'd0;
	Fy<=10'd0;
	number<=6'd0;
	is_inside<=1'b0;
	valid<=1'b0;
	 end
	else begin
	state<=next_state;
	Tx<=nTx;
	Ty<=nTy;
	Ax<=nAx;
	Ay<=nAy;
	Bx<=nBx;
	By<=nBy;
	Cx<=nCx;
	Cy<=nCy;
	Dx<=nDx;
	Dy<=nDy;
	Ex<=nEx;
	Ey<=nEy;
	Fx<=nFx;
	Fy<=nFy;
	number<=nnumber;
	is_inside<=n_inside;
	valid<=n_valid;
	end
always@(*)begin
	case(state)
		S0:begin
			next_state=S1;
			nTx=X;
			nTy=Y;
			nAx=10'd0;
			nAy=10'd0;
			nBx=10'd0;
			nBy=10'd0;
			nCx=10'd0;
			nCy=10'd0;
			nDx=10'd0;
			nDy=10'd0;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=10'd0;
			Xy=10'd0;
			Yx=10'd0;
			Yy=10'd0;
			TAx=10'd0;
			TAy=10'd0;
			TBx=10'd0;
			TBy=10'd0;
			nnumber=6'd0;
	   end
	   
		S1:begin
			nTx=Tx;
			nTy=Ty;
			nAx=X;
			nAy=Y;
			nBx=10'd0;
			nBy=10'd0;
			nCx=10'd0;
			nCy=10'd0;
			nDx=10'd0;
			nDy=10'd0;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=10'd0;
			Xy=10'd0;
			Yx=10'd0;
			Yy=10'd0;
			TAx=10'd0;
			TAy=10'd0;
			TBx=10'd0;
			TBy=10'd0;
			nnumber=6'd0;
			next_state=S2;
		end
	   
		S2:begin 
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=X;
			nBy=Y;
			nCx=10'd0;
			nCy=10'd0;
			nDx=10'd0;
			nDy=10'd0;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=10'd0;
			Xy=10'd0;
			Yx=10'd0;
			Yy=10'd0;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			next_state=S3;
		end
	   
		S3:begin 
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=X;
			nCy=Y;
			nDx=10'd0;
			nDy=10'd0;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			next_state=S4;
		end
		
		S4:begin 
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=(IO)?Bx:Cx;
			nBy=(IO)?By:Cy;
			nCx=(IO)?Cx:Bx;
			nCy=(IO)?Cy:By;
			nDx=X;
			nDy=Y;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			next_state=S5;
		end
		
		S5:begin 
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=(IO)?Cx:Dx;
			nCy=(IO)?Cy:Dy;
			nDx=(IO)?Dx:Cx;
			nDy=(IO)?Dy:Cy;
			nEx=X;
			nEy=Y;
			nFx=10'd0;
			nFy=10'd0;
			Xx=Cx;
			Xy=Cy;
			Yx=Dx;
			Yy=Dy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			next_state=S6;
		end
	
		S6:begin 
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=(IO)?Dx:Ex;
			nDy=(IO)?Dy:Ey;
			nEx=(IO)?Ex:Dx;
			nEy=(IO)?Ey:Dy;
			nFx=X;
			nFy=Y;
			Xx=Dx;
			Xy=Dy;
			Yx=Ex;
			Yy=Ey;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			next_state=5'd11;
		end
		5'd11:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nDx=Dx;
			nDy=Dy;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Ex;
			Xy=Ey;
			Yx=Fx;
			Yy=Fy;
			next_state=5'd12;
			nEx=(IO)?Ex:Fx;
			nEy=(IO)?Ey:Fy;
			nFx=(IO)?Fx:Ex;
			nFy=(IO)?Fy:Ey;
			end
		5'd12:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			nDx=Dx;
			nDy=Dy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			next_state=5'd13;
			nBx=(IO)?Bx:Cx;
			nBy=(IO)?By:Cy;
			nCx=(IO)?Cx:Bx;
			nCy=(IO)?Cy:By;
			end
		5'd13:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Cx;
			Xy=Cy;
			Yx=Dx;
			Yy=Dy;
			next_state=5'd14;
			nCx=(IO)?Cx:Dx;
			nCy=(IO)?Cy:Dy;
			nDx=(IO)?Dx:Cx;
			nDy=(IO)?Dy:Cy;
			end
		5'd14:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nFx=Fx;
			nFy=Fy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Dx;
			Xy=Dy;
			Yx=Ex;
			Yy=Ey;
			next_state=5'd15;
			nDx=(IO)?Dx:Ex;
			nDy=(IO)?Dy:Ey;
			nEx=(IO)?Ex:Dx;
			nEy=(IO)?Ey:Dy;
			end
		5'd15:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			nDx=Dx;
			nDy=Dy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			next_state=5'd16;
			nBx=(IO)?Bx:Cx;
			nBy=(IO)?By:Cy;
			nCx=(IO)?Cx:Bx;
			nCy=(IO)?Cy:By;
			end
		5'd16:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Cx;
			Xy=Cy;
			Yx=Dx;
			Yy=Dy;
			next_state=5'd17;
			nCx=(IO)?Cx:Dx;
			nCy=(IO)?Cy:Dy;
			nDx=(IO)?Dx:Cx;
			nDy=(IO)?Dy:Cy;
			end
		5'd17:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			nDx=Dx;
			nDy=Dy;
			TAx=Ax;
			TAy=Ay;
			TBx=Ax;
			TBy=Ay;
			nnumber=6'd0;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			next_state=5'd18;
			nBx=(IO)?Bx:Cx;
			nBy=(IO)?By:Cy;
			nCx=(IO)?Cx:Bx;
			nCy=(IO)?Cy:By;
			end
		5'd18:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			Xx=Ax;
			Xy=Ay;
			Yx=Bx;
			Yy=By;
			next_state=5'd19;
			nnumber[0]=IO;
			nnumber[5:1]=number[5:1];
			TAx=Tx;
			TAy=Ty;
			TBx=Ax;
			TBy=Ay;
			end
		5'd19:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Bx;
			Xy=By;
			Yx=Cx;
			Yy=Cy;
			next_state=5'd20;
			nnumber[1]=IO;
			nnumber[5:2]=number[5:2];
			nnumber[0]=number[0];
			TBx=Bx;
			TBy=By;
			end
		5'd20:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Cx;
			Xy=Cy;
			Yx=Dx;
			Yy=Dy;
			next_state=5'd21;
			nnumber[2]=IO;
			nnumber[5:3]=number[5:3];
			nnumber[1:0]=number[1:0];
			TBx=Cx;
			TBy=Cy;
			end
		5'd21:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Dx;
			Xy=Dy;
			Yx=Ex;
			Yy=Ey;
			next_state=5'd22;
			nnumber[3]=IO;
			nnumber[2:0]=number[2:0];
			nnumber[5:4]=number[5:4];
			TBx=Dx;
			TBy=Dy;
			end
		5'd22:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Ex;
			Xy=Ey;
			Yx=Fx;
			Yy=Fy;
			next_state=5'd23;
			nnumber[4]=IO;
			nnumber[3:0]=number[3:0];
			nnumber[5]=number[5];
			TBx=Ex;
			TBy=Ey;
			end
		5'd23:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Fx;
			Xy=Fy;
			Yx=Ax;
			Yy=Ay;
			next_state=5'd24;
			nnumber[5]=IO;
			nnumber[4:0]=number[4:0];
			TBx=Fx;
			TBy=Fy;
			end
		5'd24:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=Fx;
			Xy=Fy;
			Yx=Ax;
			Yy=Ay;
			next_state=5'd25;
			nnumber=number;
			TBx=Fx;
			TBy=Fy;
			end
		5'd25:begin
			nTx=Tx;
			nTy=Ty;
			nAx=Ax;
			nAy=Ay;
			nBx=Bx;
			nBy=By;
			nCx=Cx;
			nCy=Cy;
			nDx=Dx;
			nDy=Dy;
			nEx=Ex;
			nEy=Ey;
			nFx=Fx;
			nFy=Fy;
			TAx=Tx;
			TAy=Ty;
			Xx=10'd0;
			Xy=10'd0;
			Yx=10'd0;
			Yy=10'd0;
			TAx=10'd0;
			TAy=10'd0;
			TBx=10'd0;
			TBy=10'd0;
			nnumber=6'd0;
			next_state=5'd0;
			end
		default:begin
			nTx=Tx;
			nTy=Ty;
			nAx=10'd0;
			nAy=10'd0;
			nBx=10'd0;
			nBy=10'd0;
			nCx=10'd0;
			nCy=10'd0;
			nDx=10'd0;
			nDy=10'd0;
			nEx=10'd0;
			nEy=10'd0;
			nFx=10'd0;
			nFy=10'd0;
			Xx=10'd0;
			Xy=10'd0;
			Yx=10'd0;
			Yy=10'd0;
			TAx=10'd0;
			TAy=10'd0;
			TBx=10'd0;
			TBy=10'd0;
			nnumber=6'd0;
			next_state=S0;
			end
		endcase
end

endmodule